//Write a constraint for 4-bit dyanamic array. The size of the array should be in between 15 to 20.
// There should be even number in odd locations and odd number in even locations.
